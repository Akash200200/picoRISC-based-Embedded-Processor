//-----------------------------------------------------
// File Name : alucodes.sv
// Author: Akash Biyani
// Last rev. 19 Apr 2024
//-----------------------------------------------------

`define RA 3'b000
`define RB 3'b001
`define RADD 3'b010
`define RSUB 3'b011
`define RMUL 3'b100
`define RNOP 3'b101
